library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use WORK.CPU_PKG.ALL;

-- This file implements a Load-Store Unit with Total Store Ordering(TSO).
-- Store instructions are executed in-order and only after they are retired.
-- Load instructions also happen in-order but don't need to retire beforehand.

entity load_store_unit_to is
    port(
        uop_in : in T_uop;
        uop_out : out T_uop;
        cdb : in T_uop;

        agu_port : in T_lsu_gen_port;

        bus_req : out T_bus_request;
        bus_resp : in T_bus_response;
        bus_ready : in std_logic;

        stall_in : in std_logic;
        stall_out : out std_logic;

        clk : in std_logic;
        reset : in std_logic
    );
end load_store_unit_to;

architecture rtl of load_store_unit_to is
    type T_store_queue is array (0 to SQ_ENTRIES - 1) of T_lsu_store;
    signal M_store_queue : T_store_queue;
    type T_load_queue is array (0 to LQ_ENTRIES - 1) of T_lsu_load;
    signal M_load_queue : T_load_queue;

    -- STORE QUEUE CONTROL SIGNALS
    signal R_sq_head : unsigned(SQ_TAG_WIDTH - 1 downto 0);
    signal R_sq_tail : unsigned(SQ_TAG_WIDTH - 1 downto 0);
    signal R_sq_util : unsigned(SQ_TAG_WIDTH downto 0);
    signal sq_head_next : unsigned(SQ_TAG_WIDTH - 1 downto 0);
    signal sq_tail_next : unsigned(SQ_TAG_WIDTH - 1 downto 0);
    signal sq_util_next : unsigned(SQ_TAG_WIDTH downto 0);

    signal sq_head_uop : T_lsu_store;
    signal sq_head_dispatch_enable : std_logic;

    signal sq_full : std_logic;
    signal sq_empty : std_logic;

    signal sq_enqueue : std_logic;
    signal sq_dequeue : std_logic;
begin
    sq_enqueue <= not sq_full and uop_in.valid;
    sq_dequeue <= not sq_empty and sq_head_uop.retired and sq_head_uop.done;

    P_sq_next_calc : process(R_sq_head, R_sq_tail, R_sq_util, sq_enqueue, sq_dequeue)
    begin
        if R_sq_head = SQ_ENTRIES - 1 then
            sq_head_next <= (others => '0');
        else
            sq_head_next <= R_sq_head + 1;
        end if;

        if R_sq_tail = SQ_ENTRIES - 1 then
            sq_tail_next <= (others => '0');
        else
            sq_tail_next <= R_sq_tail + 1;
        end if;

        if sq_enqueue = '1' and sq_dequeue = '0' then
            sq_util_next <= R_sq_util + 1;
        elsif sq_enqueue = '0' and sq_dequeue = '1' then
            sq_util_next <= R_sq_util - 1;
        else
            sq_util_next <= R_sq_util;
        end if;
    end process;

    P_sq_cntrl : process(clk)
    begin
        if rising_edge(clk) then
            if reset = '1' then
                R_sq_head <= (others => '0');
                R_sq_tail <= (others => '0');
                R_sq_util <= (others => '0');
            else
                if agu_port.is_store = '1' then
                    -- Once the address is generated by the AGU put it into the SQ
                    if agu_port.address_valid = '1' then
                        M_store_queue(to_integer(agu_port.sq_tag)).address <= agu_port.address;
                        M_store_queue(to_integer(agu_port.sq_tag)).address_valid <= '1';
                    end if;
                    -- Once the data is generated by the AGU put it into the SQ
                    if agu_port.data_valid = '1' then
                        M_store_queue(to_integer(agu_port.sq_tag)).data <= agu_port.data;
                        M_store_queue(to_integer(agu_port.sq_tag)).data_valid <= '1';
                    end if;
                end if;

                if sq_enqueue = '1' then
                    R_sq_tail <= sq_tail_next;

                    M_store_queue(to_integer(R_sq_tail)).address <= (others => '0');
                    M_store_queue(to_integer(R_sq_tail)).address_valid <= '0';
                    M_store_queue(to_integer(R_sq_tail)).data <= (others => '0');
                    M_store_queue(to_integer(R_sq_tail)).data_valid <= '0';
                    M_store_queue(to_integer(R_sq_tail)).dispatched <= '0';
                    M_store_queue(to_integer(R_sq_tail)).done <= '0';
                    M_store_queue(to_integer(R_sq_tail)).retired <= '1';
                end if;
                
                if bus_ready = '1' and sq_head_dispatch_enable = '1' then
                    M_store_queue(to_integer(R_sq_head)).dispatched <= '1';
                end if;

                if bus_resp.valid = '1' then
                    M_store_queue(to_integer(R_sq_head)).done <= '1';
                end if;

                if sq_dequeue = '1' then
                    R_sq_head <= sq_head_next;
                end if;

                R_sq_util <= sq_util_next;
            end if;
        end if;
    end process;
    sq_head_uop <= M_store_queue(to_integer(R_sq_head));
    sq_head_dispatch_enable <= sq_head_uop.data_valid and sq_head_uop.address_valid and not sq_head_uop.dispatched and sq_head_uop.retired;

    bus_req.address <= sq_head_uop.address;
    bus_req.data <= sq_head_uop.data;
    bus_req.data_size <= "00";
    bus_req.is_store <= '1';
    bus_req.sq_tag <= R_sq_head;
    bus_req.lq_tag <= (others => '0');
    bus_req.valid <= sq_head_dispatch_enable;

    sq_full <= '1' when R_sq_util = SQ_ENTRIES else '0';
    sq_empty <= '1' when R_sq_util = 0 else '0';

    stall_out <= sq_full;
end rtl;
