library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity cpu_core is

end cpu_core;

architecture rtl of cpu_core is

begin


end rtl;
