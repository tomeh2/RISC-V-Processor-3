library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity scheduler is

end scheduler;

architecture rtl of scheduler is

begin

end rtl;
