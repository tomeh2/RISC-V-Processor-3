library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity execution_unit is

end execution_unit;

architecture rtl of execution_unit is

begin

end rtl;
