library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity front_end is

end front_end;

architecture rtl of front_end is

begin


end rtl;
