library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity back_end is

end back_end;

architecture rtl of back_end is

begin


end rtl;
