library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity cpu is

end cpu;

architecture rtl of cpu is

begin


end rtl;
