library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity top_sim is

end top_sim;

architecture Behavioral of top_sim is

begin


end Behavioral;
