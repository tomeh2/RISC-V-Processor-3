library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package cpu_pkg is
    
end package;
